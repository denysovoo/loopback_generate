library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;

entity bram_tdp is
generic (
    DATA    : integer := 32;
    ADDR    : integer := 8
);
port (
    -- Port A
    a_clk   : in  std_logic;
    a_wr    : in  std_logic;
    a_addr  : in  std_logic_vector(ADDR-1 downto 0);
    a_din   : in  std_logic_vector(DATA-1 downto 0);
    a_dout  : out std_logic_vector(DATA-1 downto 0);

    -- Port B
    b_clk   : in  std_logic;
    b_wr    : in  std_logic;
    b_addr  : in  std_logic_vector(ADDR-1 downto 0);
    b_din   : in  std_logic_vector(DATA-1 downto 0);
    b_dout  : out std_logic_vector(DATA-1 downto 0)
);
end bram_tdp;

architecture rtl of bram_tdp is
    -- Shared memory
    type mem_type is array ( (2**ADDR)-1 downto 0 ) of std_logic_vector(DATA-1 downto 0);
    
   -- FUNCTION initialize_ram  return mem_type is variable result : mem_type;
   -- BEGIN
		-- FOR i IN ((2**ADDR)-1) DOWNTO 0 LOOP
			-- result(i) := std_logic_vector( to_unsigned(natural(i), natural'(DATA)));
		-- END LOOP;
   -- RETURN result;
   -- END initialize_ram;
	
	shared variable mem : mem_type;
    
--    shared variable mem : mem_type := 
--(	--"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	"00000000000000000000000000000000",
--	
--	"00000000000000000000000000001101",
--	"00000000000000000000000011110011",--
--	"00000000000000000000000000000101",
--	"00000000000000000000000011110000",--
--	"00000000000000000000000000000111",
--	"00000000000000000000000010110000",--
--	"00000000000000000000000000000011",
--	"00000000000000000000000010010000",--
--
--	"00000000000000000000000000000101",
--	"00000000000000000000000011110000",--
--	"00000000000000000000000000000111",
--	"00000000000000000000000010110000",--
--	"00000000000000000000000000000011",
--	"00000000000000000000000010010000",--
--	
--	"00000000000000000000000000001000", --add now!!! -- it's normal speed
--	
--	"00000000000000000000011111111111",
--	"00000000000000000000000000010000",
--	"00000000000000000000000000000011",
--	"00000000000000000000000000000011"
--	
--	); -- := initialize_ram; --mem_type

	begin

-- Port A
process(a_clk)
begin
    if(a_clk'event and a_clk='1') then
        if(a_wr='1') then
            mem(conv_integer(a_addr)) := a_din;
        end if;
        a_dout <= mem(conv_integer(a_addr));
    end if;
end process;

-- Port B
process(b_clk)
begin
    if(b_clk'event and b_clk='1') then
        if(b_wr='1') then
            mem(conv_integer(b_addr)) := b_din;
        end if;
        b_dout <= mem(conv_integer(b_addr));
    end if;
end process;

end rtl;